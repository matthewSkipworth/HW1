module Mux_5_to_1(S, U, V, W, X, Y, M);
	input U, V, W, X, Y;
	input [2:0] S;
	output reg M;
	
	wire A, B, C;
	//module Mux_2_to_1(S, X, Y, M);
/*	Mux_2_to_1 M0(S[0], U, V, A);
	Mux_2_to_1 M1(S[0], W, X, B);
	Mux_2_to_1 M2(S[1], A, B, C);
	Mux_2_to_1 M3(S[2], C, Y, M);*/
	assign A = (~S[0] & U) | (S[0] & V);
	assign B = (~S[0] & W) | (S[0] & X);
	assign C = (~S[1] & A) | (S[1] & B);
	assign M = (~S[2] & C) | (S[2] & Y);
endmodule

//module Mux_5_to_1_testbench(input  U, V, W, X, Y, [2:0] S,output reg M);
module Mux_5_to_1_testbench();
	logic U;
	logic V;
	logic W; 
	logic X;
	logic Y; 
	logic M;
	logic [2:0] S;
	Mux_5_to_1 dut(.S(S), .U(U), .V(V), .W(W), .X(X), .Y(Y), .M(M));
	initial begin
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 0; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 0; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 0; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 0; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 0; W = 1; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 0; X = 1; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 0; Y = 1; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 0; M = 1; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 0; #10;
	S[0] = 1; S[1] = 1; S[2] = 1; U = 1; V = 1; W = 1; X = 1; Y = 1; M = 1; #10;
	end
endmodule